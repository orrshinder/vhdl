-- megafunction wizard: %PLL Intel FPGA IP v20.1%
-- GENERATION: XML
-- clock_generator.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity clock_generator is
	port (
		refclk   : in  std_logic := '0'; --  refclk.clk
		rst      : in  std_logic := '0'; --   reset.reset
		outclk_0 : out std_logic;        -- outclk0.clk
		locked   : out std_logic         --  locked.export
	);
end entity clock_generator;

architecture rtl of clock_generator is

	constant C_CLK_PRD	: time := 40 ns;

	signal clk_sig		: std_logic := 'X';
	signal locked_int	: std_logic := '0';

begin	
	
	process
	begin
	
		locked_int <= '0';
		wait until rst = '0';
		wait for 10 us;
		locked_int <= '1';
		wait until rst = '0';
		
	end process;

	process
	begin
		wait until locked_int = '1';
		
		while locked_int = '1' loop
			clk_sig <= '1';
			wait for C_CLK_PRD / 2;
			clk_sig <= '0';
			wait for C_CLK_PRD / 2;
		end loop;
		
		clk_sig <= 'X';
	end process;
	
	outclk_0 <= clk_sig;
	
	process
	begin
		locked <= '0';
		wait until locked_int  = '1';
		wait for 100 ns;
		wait until rising_edge(clk_sig);
		locked <= '1';
		wait until locked_int = '0';
		locked <= '0';
	end process;
		
end architecture;